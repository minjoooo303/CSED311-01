`include "opcodes.v"

module immediate_generator (    input [31:0] instr,
                                output reg [31:0] imm_gen_out );

    always @(*) begin //조합논리 블록이므로 블로킹 할당 사용
        case(instr[6:0])
            `ARITHMETIC: begin // R-type
                imm_gen_out = 32'b0;
            end
            `ARITHMETIC_IMM, `LOAD, `JALR: begin // I-type
                imm_gen_out = {{20{instr[31]}}, instr[31:20]}; //부호 확장을 함
            end
            `STORE: begin // S-type
                imm_gen_out = {{20{instr[31]}}, instr[31:25], instr[11:7]};
            end
            `BRANCH: begin // SB-type
                imm_gen_out = {{19{inst[31]}}, instr[31], instr[7], instr[30:25], instr[11:8], 1'b0}
            end
            `JAL: begin // J-type
                imm_gen_out = {{11{instr[31]}}, instr[31], instr[19:12], instr[20], instr[30:21], 1'b0}
            end
            default: begin
                imm_gen_out = 32'b0;
            end

        endcase
    end


endmodule